library verilog;
use verilog.vl_types.all;
entity reciprocal_tbb is
end reciprocal_tbb;
