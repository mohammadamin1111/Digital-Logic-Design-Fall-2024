module multiplier(input signed [7:0] x,input signed [7:0] y,output signed [15:0] multiplier_result);
       assign multiplier_result =x*y;
endmodule
