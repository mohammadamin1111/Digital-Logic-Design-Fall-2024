module one_hot_encoder(input [15:0] w, output reg signed [3:0] y);

  always @(*) 
    begin
      case (w)
        16'b1000000000000000: y = -8;
        16'b0100000000000000: y = -7;
        16'b0010000000000000: y = -6;
        16'b0001000000000000: y = -5;
        16'b0000100000000000: y = -4;
        16'b0000010000000000: y = -3;
        16'b0000001000000000: y = -2;
        16'b0000000100000000: y = -1;
        16'b0000000010000000: y = 0;
        16'b0000000001000000: y = 1;
        16'b0000000000100000: y = 2;
        16'b0000000000010000: y = 3;
        16'b0000000000001000: y = 4;
        16'b0000000000000100: y = 5;
        16'b0000000000000010: y = 6;
        16'b0000000000000001: y = 7;
        
      endcase
    end
endmodule
